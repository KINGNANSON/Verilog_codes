

module helloworld();

initial begin
    $display("Hello I am Nanson , course start date is 27 JUne 2023");
end

endmodule
